module log

pub const false_log := '\033[31m[False] \033[0m'
pub const true_log := '\033[32m[True] \033[0m'
pub const warn_log := '\033[33m[Warn] \033[0m'



