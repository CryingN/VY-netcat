module client

pub struct SetServer {
pub:
	exec		string
	security	string
pub mut:
	port		string
	keep		bool
}

